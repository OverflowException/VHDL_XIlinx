----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:17:53 11/08/2017 
-- Design Name: 
-- Module Name:    display - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity display_tkr is
	port(
			number: in std_logic_vector(3 downto 0);
			segs: out std_logic_vector(7 downto 0));
end display_tkr;

architecture Behavioral of display_tkr is 
begin
    with number Select
		segs(7 downto 0) <= 
			"11000000" when "0000",   --0
			"11111001" when "0001",   --1
         "10100100" when "0010",   --2
         "10110000" when "0011",   --3
         "10011001" when "0100",   --4
         "10010010" when "0101",   --5
         "10000010" when "0110",   --6
         "11111000" when "0111",   --7
         "10000000" when "1000",   --8
         "10010000" when "1001",   --9
         "10001000" when "1010",   --A
         "10000011" when "1011",   --b
         "10000111" when "1100",   --t(C)
         "10001001" when "1101",   --K(D)
         "10000110" when "1110",   --E(E)
         "10101111" when "1111",   --r(F)
         "11000000" when others;   --0
			
end Behavioral;

